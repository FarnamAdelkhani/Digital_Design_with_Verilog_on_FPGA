library verilog;
use verilog.vl_types.all;
entity testArith is
end testArith;
