library verilog;
use verilog.vl_types.all;
entity Testbench_1 is
end Testbench_1;
