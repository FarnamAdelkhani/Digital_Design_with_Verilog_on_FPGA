library verilog;
use verilog.vl_types.all;
entity testDlatch is
end testDlatch;
