library verilog;
use verilog.vl_types.all;
entity bitTest is
end bitTest;
