library verilog;
use verilog.vl_types.all;
entity TestArith is
end TestArith;
