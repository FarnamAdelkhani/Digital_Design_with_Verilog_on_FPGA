library verilog;
use verilog.vl_types.all;
entity testJK is
end testJK;
